LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

LIBRARY STD;
USE STD.ALL;

ENTITY bsim3_addnoise IS
  GENERIC (
   w :   real :=  5.000000e-06;
   l :   real :=  5.000000e-06;
   \_m\ :   real :=  1.000000e+00;
   paramchk :   integer  := 1;
   PMOS :   integer  := 0;
   vth0 :   real :=  -9.999900e-99;
   vfb :   real :=  -9.999900e-99;
   k1 :   real :=  -9.999900e-99;
   k2 :   real :=  -9.999900e-99;
   k3 :   integer  := 80;
   k3b :   integer  := 0;
   w0 :   real :=  2.500000e-06;
   nlx :   real :=  1.740000e-07;
   gamma1 :   real :=  -9.999900e-99;
   gamma2 :   real :=  0.000000e+00;
   vbx :   real :=  -9.999900e-99;
   vbm :   integer  := -3;
   dvt0 :   real :=  2.200000e+00;
   dvt1 :   real :=  5.300000e-01;
   dvt2 :   real :=  -3.200000e-02;
   dvt0w :   integer  := 0;
   dvt1w :   real :=  5.300000e+06;
   dvt2w :   real :=  -3.200000e-02;
   a0 :   integer  := 1;
   b0 :   integer  := 0;
   b1 :   integer  := 0;
   a1 :   integer  := 0;
   a2 :   integer  := 1;
   ags :   integer  := 0;
   keta :   real :=  -4.700000e-02;
   nsub :   real :=  -9.999900e-99;
   nch :   real :=  -9.999900e-99;
   ngate :   real :=  -9.999900e-99;
   xj :   real :=  1.500000e-07;
   lint :   integer  := 0;
   wint :   integer  := 0;
   ll :   integer  := 0;
   lln :   integer  := 1;
   lw :   integer  := 0;
   lwn :   integer  := 1;
   lwl :   integer  := 0;
   wl :   integer  := 0;
   wln :   integer  := 1;
   ww :   integer  := 0;
   wwn :   integer  := 1;
   wwl :   integer  := 0;
   dwg :   integer  := 0;
   dwb :   integer  := 0;
   tox :   real :=  1.500000e-08;
   xt :   real :=  -9.999900e-99;
   rdsw :   integer  := 0;
   prwb :   integer  := 0;
   prwg :   integer  := 0;
   wr :   integer  := 1;
   binunit :   integer  := 1;
   mobmod :   integer  := 1;
   u0 :   real :=  -9.999900e-99;
   vsat :   real :=  8.000000e+04;
   ua :   real :=  2.250000e-09;
   ub :   real :=  5.870000e-19;
   uc :   real :=  -9.999900e-99;
   drout :   real :=  5.600000e-01;
   pclm :   real :=  1.300000e+00;
   pdiblc1 :   real :=  3.900000e-01;
   pdiblc2 :   real :=  8.600000e-03;
   pdiblcb :   real :=  0.000000e+00;
   pscbe1 :   real :=  4.240000e+08;
   pscbe2 :   real :=  1.000000e-05;
   pvag :   integer  := 0;
   delta :   real :=  1.000000e-02;
   cdsc :   real :=  2.400000e-04;
   cdscb :   integer  := 0;
   cdscd :   integer  := 0;
   nfactor :   integer  := 1;
   cit :   integer  := 0;
   voff :   real :=  -8.000000e-02;
   eta0 :   real :=  8.000000e-02;
   etab :   real :=  -7.000000e-02;
   xpart :   integer  := 0;
   capmod :   integer  := 3;
   dlc :   real :=  -9.999900e-99;
   clc :   real :=  1.000000e-07;
   cle :   real :=  6.000000e-01;
   vfbcv :   integer  := -1;
   acde :   integer  := 1;
   moin :   integer  := 15;
   noff :   integer  := 1;
   voffcv :   integer  := 0;
   tnom :   integer  := 27;
   kt1 :   real :=  -1.100000e-01;
   kt1l :   integer  := 0;
   kt2 :   real :=  2.200000e-02;
   at :   real :=  3.300000e+04;
   ua1 :   real :=  4.310000e-09;
   ub1 :   real :=  -7.610000e-18;
   uc1 :   real :=  -9.999900e-99;
   prt :   integer  := 0;
   ute :   real :=  -1.500000e+00;
   noimod :   integer  := 1;
   ntnoi :   real :=  1.000000e+00;
   dlclm :   real :=  0.000000e+00;
   wmax :   integer  := 1;
   wmin :   integer  := 0;
   lmax :   integer  := 1;
   lmin :   integer  := 0;
   xl :   integer  := 0;
   xw :   integer  := 0;
   lcdsc :   real :=  0.000000e+00;
   lcdscb :   real :=  0.000000e+00;
   lcdscd :   real :=  0.000000e+00;
   lcit :   real :=  0.000000e+00;
   lnfactor :   real :=  0.000000e+00;
   lxj :   real :=  0.000000e+00;
   lvsat :   real :=  0.000000e+00;
   lat :   real :=  0.000000e+00;
   la0 :   real :=  0.000000e+00;
   lags :   real :=  0.000000e+00;
   la1 :   real :=  0.000000e+00;
   la2 :   real :=  0.000000e+00;
   lketa :   real :=  0.000000e+00;
   lnsub :   real :=  0.000000e+00;
   lnch :   real :=  0.000000e+00;
   lngate :   real :=  0.000000e+00;
   lgamma1 :   real :=  0.000000e+00;
   lgamma2 :   real :=  0.000000e+00;
   lvbx :   real :=  0.000000e+00;
   lvbm :   real :=  0.000000e+00;
   lxt :   real :=  0.000000e+00;
   lk1 :   real :=  0.000000e+00;
   lkt1 :   real :=  0.000000e+00;
   lkt1l :   real :=  0.000000e+00;
   lkt2 :   real :=  0.000000e+00;
   lk2 :   real :=  0.000000e+00;
   lk3 :   real :=  0.000000e+00;
   lk3b :   real :=  0.000000e+00;
   lw0 :   real :=  0.000000e+00;
   lnlx :   real :=  0.000000e+00;
   ldvt0 :   real :=  0.000000e+00;
   ldvt1 :   real :=  0.000000e+00;
   ldvt2 :   real :=  0.000000e+00;
   ldvt0w :   real :=  0.000000e+00;
   ldvt1w :   real :=  0.000000e+00;
   ldvt2w :   real :=  0.000000e+00;
   ldrout :   real :=  0.000000e+00;
   ldsub :   real :=  0.000000e+00;
   lvth0 :   real :=  0.000000e+00;
   lua :   real :=  0.000000e+00;
   lua1 :   real :=  0.000000e+00;
   lub :   real :=  0.000000e+00;
   lub1 :   real :=  0.000000e+00;
   luc :   real :=  0.000000e+00;
   luc1 :   real :=  0.000000e+00;
   lu0 :   real :=  0.000000e+00;
   lute :   real :=  0.000000e+00;
   lvoff :   real :=  0.000000e+00;
   ldelta :   real :=  0.000000e+00;
   lrdsw :   real :=  0.000000e+00;
   lprwg :   real :=  0.000000e+00;
   lprwb :   real :=  0.000000e+00;
   lprt :   real :=  0.000000e+00;
   leta0 :   real :=  0.000000e+00;
   letab :   real :=  0.000000e+00;
   lpclm :   real :=  0.000000e+00;
   lpdiblc1 :   real :=  0.000000e+00;
   lpdiblc2 :   real :=  0.000000e+00;
   lpdiblcb :   real :=  0.000000e+00;
   lpscbe1 :   real :=  0.000000e+00;
   lpscbe2 :   integer  := 0;
   lpvag :   real :=  0.000000e+00;
   lwr :   real :=  0.000000e+00;
   ldwg :   real :=  0.000000e+00;
   ldwb :   real :=  0.000000e+00;
   lb0 :   real :=  0.000000e+00;
   lb1 :   real :=  0.000000e+00;
   lclc :   real :=  0.000000e+00;
   lcle :   real :=  0.000000e+00;
   lvfbcv :   real :=  0.000000e+00;
   lvfb :   real :=  0.000000e+00;
   lacde :   real :=  0.000000e+00;
   lmoin :   real :=  0.000000e+00;
   lnoff :   real :=  0.000000e+00;
   lvoffcv :   real :=  0.000000e+00;
   wcdsc :   real :=  0.000000e+00;
   wcdscb :   real :=  0.000000e+00;
   wcdscd :   real :=  0.000000e+00;
   wcit :   real :=  0.000000e+00;
   wnfactor :   real :=  0.000000e+00;
   wxj :   real :=  0.000000e+00;
   wvsat :   real :=  0.000000e+00;
   wat :   real :=  0.000000e+00;
   wa0 :   real :=  0.000000e+00;
   wags :   real :=  0.000000e+00;
   wa1 :   real :=  0.000000e+00;
   wa2 :   real :=  0.000000e+00;
   wketa :   real :=  0.000000e+00;
   wnsub :   real :=  0.000000e+00;
   wnch :   real :=  0.000000e+00;
   wngate :   real :=  0.000000e+00;
   wgamma1 :   real :=  0.000000e+00;
   wgamma2 :   real :=  0.000000e+00;
   wvbx :   real :=  0.000000e+00;
   wvbm :   real :=  0.000000e+00;
   wxt :   real :=  0.000000e+00;
   wk1 :   real :=  0.000000e+00;
   wkt1 :   real :=  0.000000e+00;
   wkt1l :   real :=  0.000000e+00;
   wkt2 :   real :=  0.000000e+00;
   wk2 :   real :=  0.000000e+00;
   wk3 :   real :=  0.000000e+00;
   wk3b :   real :=  0.000000e+00;
   ww0 :   real :=  0.000000e+00;
   wnlx :   real :=  0.000000e+00;
   wdvt0 :   real :=  0.000000e+00;
   wdvt1 :   real :=  0.000000e+00;
   wdvt2 :   real :=  0.000000e+00;
   wdvt0w :   real :=  0.000000e+00;
   wdvt1w :   real :=  0.000000e+00;
   wdvt2w :   real :=  0.000000e+00;
   wdrout :   real :=  0.000000e+00;
   wdsub :   real :=  0.000000e+00;
   wvth0 :   real :=  0.000000e+00;
   wua :   real :=  0.000000e+00;
   wua1 :   real :=  0.000000e+00;
   wub :   real :=  0.000000e+00;
   wub1 :   real :=  0.000000e+00;
   wuc :   real :=  0.000000e+00;
   wuc1 :   real :=  0.000000e+00;
   wu0 :   real :=  0.000000e+00;
   wute :   real :=  0.000000e+00;
   wvoff :   real :=  0.000000e+00;
   wdelta :   real :=  0.000000e+00;
   wrdsw :   real :=  0.000000e+00;
   wprwg :   real :=  0.000000e+00;
   wprwb :   real :=  0.000000e+00;
   wprt :   real :=  0.000000e+00;
   weta0 :   real :=  0.000000e+00;
   wetab :   real :=  0.000000e+00;
   wpclm :   real :=  0.000000e+00;
   wpdiblc1 :   real :=  0.000000e+00;
   wpdiblc2 :   real :=  0.000000e+00;
   wpdiblcb :   real :=  0.000000e+00;
   wpscbe1 :   real :=  0.000000e+00;
   wpscbe2 :   real :=  0.000000e+00;
   wpvag :   real :=  0.000000e+00;
   wwr :   real :=  0.000000e+00;
   wdwg :   real :=  0.000000e+00;
   wdwb :   real :=  0.000000e+00;
   wb0 :   real :=  0.000000e+00;
   wb1 :   real :=  0.000000e+00;
   wclc :   real :=  0.000000e+00;
   wcle :   real :=  0.000000e+00;
   wvfbcv :   real :=  0.000000e+00;
   wvfb :   real :=  0.000000e+00;
   wacde :   real :=  0.000000e+00;
   wmoin :   real :=  0.000000e+00;
   wnoff :   real :=  0.000000e+00;
   wvoffcv :   real :=  0.000000e+00;
   pcdsc :   real :=  0.000000e+00;
   pcdscb :   real :=  0.000000e+00;
   pcdscd :   real :=  0.000000e+00;
   pcit :   real :=  0.000000e+00;
   pnfactor :   real :=  0.000000e+00;
   pxj :   real :=  0.000000e+00;
   pvsat :   real :=  0.000000e+00;
   pat :   real :=  0.000000e+00;
   pa0 :   real :=  0.000000e+00;
   pags :   real :=  0.000000e+00;
   pa1 :   real :=  0.000000e+00;
   pa2 :   real :=  0.000000e+00;
   pketa :   real :=  0.000000e+00;
   pnsub :   real :=  0.000000e+00;
   pnch :   real :=  0.000000e+00;
   pngate :   real :=  0.000000e+00;
   pgamma1 :   real :=  0.000000e+00;
   pgamma2 :   real :=  0.000000e+00;
   pvbx :   real :=  0.000000e+00;
   pvbm :   real :=  0.000000e+00;
   pxt :   real :=  0.000000e+00;
   pk1 :   real :=  0.000000e+00;
   pkt1 :   real :=  0.000000e+00;
   pkt1l :   real :=  0.000000e+00;
   pkt2 :   real :=  0.000000e+00;
   pk2 :   real :=  0.000000e+00;
   pk3 :   real :=  0.000000e+00;
   pk3b :   real :=  0.000000e+00;
   pw0 :   real :=  0.000000e+00;
   pnlx :   real :=  0.000000e+00;
   pdvt0 :   real :=  0.000000e+00;
   pdvt1 :   real :=  0.000000e+00;
   pdvt2 :   real :=  0.000000e+00;
   pdvt0w :   real :=  0.000000e+00;
   pdvt1w :   real :=  0.000000e+00;
   pdvt2w :   real :=  0.000000e+00;
   pdrout :   real :=  0.000000e+00;
   pdsub :   real :=  0.000000e+00;
   pvth0 :   real :=  0.000000e+00;
   pua :   real :=  0.000000e+00;
   pua1 :   real :=  0.000000e+00;
   pub :   real :=  0.000000e+00;
   pub1 :   real :=  0.000000e+00;
   puc :   real :=  0.000000e+00;
   puc1 :   real :=  0.000000e+00;
   pu0 :   real :=  0.000000e+00;
   pute :   real :=  0.000000e+00;
   pvoff :   real :=  0.000000e+00;
   pdelta :   real :=  0.000000e+00;
   prdsw :   real :=  0.000000e+00;
   pprwg :   real :=  0.000000e+00;
   pprwb :   real :=  0.000000e+00;
   pprt :   real :=  0.000000e+00;
   peta0 :   real :=  0.000000e+00;
   petab :   real :=  0.000000e+00;
   ppclm :   real :=  0.000000e+00;
   ppdiblc1 :   real :=  0.000000e+00;
   ppdiblc2 :   real :=  0.000000e+00;
   ppdiblcb :   real :=  0.000000e+00;
   ppscbe1 :   real :=  0.000000e+00;
   ppscbe2 :   real :=  0.000000e+00;
   ppvag :   real :=  0.000000e+00;
   pwr_noise :   real :=  0.000000e+00;
   pdwg :   real :=  0.000000e+00;
   pdwb :   real :=  0.000000e+00;
   pb0 :   real :=  0.000000e+00;
   pb1 :   real :=  0.000000e+00;
   pclc :   real :=  0.000000e+00;
   pcle :   real :=  0.000000e+00;
   pvfbcv :   real :=  0.000000e+00;
   pvfb :   real :=  0.000000e+00;
   pacde :   real :=  0.000000e+00;
   pmoin :   real :=  0.000000e+00;
   pnoff :   real :=  0.000000e+00;
   pvoffcv :   real :=  0.000000e+00 );
  PORT (
    SIGNAL d : INOUT STD_LOGIC;
    SIGNAL g : INOUT STD_LOGIC;
    SIGNAL s : INOUT STD_LOGIC;
    SIGNAL b : INOUT STD_LOGIC);
END ENTITY bsim3_addnoise;

